-- ########################################################################
--! @file       link_layer_crc.vhd
--! @brief      crc generator which takes input data and outputs the calculated crc.
--! @details    Takes input data and saves intermediate crc values to compute a final crc based on a set of data.
--! @author     Hannah Mohr
--! @date       April 2017
--! @copyright  Copyright (C) 2017 Ross K. Snider and Hannah D. Mohr
--
-- CRC Engine RTL Design
-- Copyright (C) www.ElectronicDesignworks.com
-- Source code generated by ElectronicDesignworks IP Generator (CRC).
-- Documentation can be downloaded from www.ElectronicDesignworks.com
--
--  This program is free software: you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation, either version 3 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS for A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
-- ********************************
-- 			Source Code
-- ********************************
--
-- ********************************
--            License
-- ********************************
-- This source file may be used and distributed freely provided that this
-- copyright notice, list of conditions and the following disclaimer is
-- not removed from the file.
-- Any derivative work should contain this copyright notice and associated disclaimer.
-- This source code file is provided "AS IS" AND WITHOUT ANY WARRANTY,
-- without even the implied warranty of MERCHANTABILITY or FITNESS FOR A
-- PARTICULAR PURPOSE.
-- ********************************
--           Specification
-- ********************************
-- File Name       : CRC32_DATA32.vhd
-- Description     : CRC Engine ENTITY
-- Clock           : Positive Edge
-- Reset           : Active Low
-- First Serial    : MSB
-- Data Bus Width  : 32 bits
-- Polynomial      : (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
-- Date            : 18-Jan-2017
-- Version         : 1.0
-- ########################################################################

library ieee ;
use ieee.std_logic_1164.all ;
use ieee.std_logic_arith.all ;
use ieee.std_logic_unsigned.all ;

entity link_layer_crc is
   port(clk	       		: in  std_logic;
        rst_n      		: in  std_logic;
        crc_start  		: in  std_logic;									-- input signal to start the crc calculation
        crc_data_in		: in  std_logic_vector(31 downto 0);				-- input signal containing the data on which the crc is to be calculated
        crc_data_valid 	: in  std_logic;									-- input signal indicating crc_data_in is valid and the computation should proceed
        crc_out    		: out std_logic_vector(31 downto 0));				-- calculated value for the crc on the input data
end entity;

architecture behave of link_layer_crc is

 signal crc_i          	: std_logic_vector(31 downto 0);		-- initial/previous value to use in the crc calculation
 signal crc_c          	: std_logic_vector(31 downto 0);		-- output of crc calculation
 signal crc_r         	: std_logic_vector(31 downto 0);		-- output of crc calculation when input data are valid
 
 constant crc_const    	: std_logic_vector(31 downto 0) := x"52325032";		-- seed value defined by SATA protocol

begin
-- assign the value of the crc used in the calculation
crc_i    <= crc_const when crc_start = '1' else		-- initialize with the seed at start-up
            crc_r;									-- use the previously calculated crc value

-- XOR calculation to generate the crc based on the previous crc value and the input data
crc_c(0) <= crc_data_in(0) xor crc_data_in(6) xor crc_data_in(9) xor crc_data_in(10) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(28) xor crc_i(28) xor crc_i(10) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(25) xor crc_i(25) xor crc_data_in(12) xor crc_data_in(16) xor crc_data_in(30) xor crc_i(6) xor crc_i(30) xor crc_i(16) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(1) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(7) xor crc_data_in(11) xor crc_i(1) xor crc_i(11) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(13) xor crc_data_in(17) xor crc_i(7) xor crc_i(17) xor crc_i(13) xor crc_data_in(6) xor crc_data_in(9) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(28) xor crc_i(28) xor crc_i(9) xor crc_data_in(12) xor crc_data_in(16) xor crc_i(6) xor crc_i(16) xor crc_i(12);
crc_c(2) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(2) xor crc_data_in(8) xor crc_i(2) xor crc_data_in(14) xor crc_data_in(18) xor crc_i(8) xor crc_i(18) xor crc_i(14) xor crc_data_in(7) xor crc_i(1) xor crc_data_in(13) xor crc_data_in(17) xor crc_i(7) xor crc_i(17) xor crc_i(13) xor crc_data_in(6) xor crc_data_in(9) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(16) xor crc_data_in(30) xor crc_i(6) xor crc_i(30) xor crc_i(16) xor crc_data_in(31) xor crc_i(31);
crc_c(3) <= crc_data_in(1) xor crc_data_in(2) xor crc_data_in(3) xor crc_data_in(9) xor crc_i(3) xor crc_data_in(15) xor crc_data_in(19) xor crc_i(9) xor crc_i(19) xor crc_i(15) xor crc_data_in(8) xor crc_i(2) xor crc_data_in(14) xor crc_data_in(18) xor crc_i(8) xor crc_i(18) xor crc_i(14) xor crc_data_in(7) xor crc_data_in(10) xor crc_data_in(25) xor crc_i(1) xor crc_i(25) xor crc_data_in(27) xor crc_i(27) xor crc_i(10) xor crc_data_in(17) xor crc_data_in(31) xor crc_i(7) xor crc_i(31) xor crc_i(17);
crc_c(4) <= crc_data_in(0) xor crc_data_in(2) xor crc_data_in(3) xor crc_data_in(4) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_i(3) xor crc_data_in(15) xor crc_data_in(19) xor crc_i(19) xor crc_i(15) xor crc_data_in(8) xor crc_data_in(11) xor crc_i(2) xor crc_i(11) xor crc_data_in(18) xor crc_i(8) xor crc_i(18) xor crc_data_in(6) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(25) xor crc_i(25) xor crc_data_in(12) xor crc_data_in(30) xor crc_i(6) xor crc_i(30) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(5) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(3) xor crc_data_in(4) xor crc_data_in(5) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_i(3) xor crc_data_in(19) xor crc_i(19) xor crc_data_in(7) xor crc_i(1) xor crc_data_in(13) xor crc_i(7) xor crc_i(13) xor crc_data_in(6) xor crc_data_in(10) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(28) xor crc_i(28) xor crc_i(10) xor crc_i(6);
crc_c(6) <= crc_data_in(1) xor crc_data_in(2) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(6) xor crc_i(6) xor crc_data_in(22) xor crc_i(22) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_data_in(8) xor crc_i(2) xor crc_data_in(14) xor crc_i(8) xor crc_i(14) xor crc_data_in(7) xor crc_data_in(11) xor crc_data_in(25) xor crc_i(1) xor crc_i(25) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(29) xor crc_i(29) xor crc_i(11) xor crc_i(7);
crc_c(7) <= crc_data_in(0) xor crc_data_in(2) xor crc_data_in(3) xor crc_data_in(5) xor crc_data_in(7) xor crc_i(7) xor crc_data_in(23) xor crc_i(23) xor crc_data_in(22) xor crc_i(22) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_i(3) xor crc_data_in(15) xor crc_i(15) xor crc_data_in(8) xor crc_i(2) xor crc_i(8) xor crc_data_in(10) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(28) xor crc_i(28) xor crc_i(10) xor crc_data_in(25) xor crc_i(25) xor crc_data_in(16) xor crc_i(16);
crc_c(8) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(3) xor crc_data_in(4) xor crc_data_in(8) xor crc_i(8) xor crc_data_in(23) xor crc_i(23) xor crc_data_in(22) xor crc_i(22) xor crc_i(4) xor crc_i(3) xor crc_data_in(11) xor crc_i(1) xor crc_i(11) xor crc_data_in(17) xor crc_i(17) xor crc_data_in(10) xor crc_i(0) xor crc_data_in(28) xor crc_i(28) xor crc_i(10) xor crc_data_in(12) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(9) <= crc_data_in(1) xor crc_data_in(2) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(9) xor crc_i(9) xor crc_data_in(24) xor crc_i(24) xor crc_data_in(23) xor crc_i(23) xor crc_i(5) xor crc_i(4) xor crc_data_in(12) xor crc_i(2) xor crc_i(12) xor crc_data_in(18) xor crc_i(18) xor crc_data_in(11) xor crc_i(1) xor crc_data_in(29) xor crc_i(29) xor crc_i(11) xor crc_data_in(13) xor crc_i(13);
crc_c(10) <= crc_data_in(0) xor crc_data_in(2) xor crc_data_in(3) xor crc_data_in(5) xor crc_i(5) xor crc_data_in(13) xor crc_i(3) xor crc_i(13) xor crc_data_in(19) xor crc_i(19) xor crc_i(2) xor crc_data_in(14) xor crc_i(14) xor crc_data_in(9) xor crc_i(0) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(16) xor crc_i(16) xor crc_data_in(31) xor crc_i(31);
crc_c(11) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(3) xor crc_data_in(4) xor crc_data_in(14) xor crc_i(4) xor crc_i(14) xor crc_data_in(20) xor crc_i(20) xor crc_i(3) xor crc_data_in(15) xor crc_i(15) xor crc_i(1) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(17) xor crc_i(17) xor crc_data_in(9) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(25) xor crc_i(25) xor crc_data_in(12) xor crc_data_in(16) xor crc_i(16) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(12) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(2) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(15) xor crc_i(5) xor crc_i(15) xor crc_data_in(21) xor crc_i(21) xor crc_i(4) xor crc_i(2) xor crc_data_in(18) xor crc_i(18) xor crc_i(1) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(13) xor crc_data_in(17) xor crc_i(17) xor crc_i(13) xor crc_data_in(6) xor crc_data_in(9) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_i(9) xor crc_data_in(12) xor crc_data_in(30) xor crc_i(6) xor crc_i(30) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(13) <= crc_data_in(1) xor crc_data_in(2) xor crc_data_in(3) xor crc_data_in(5) xor crc_data_in(6) xor crc_data_in(16) xor crc_i(6) xor crc_i(16) xor crc_data_in(22) xor crc_i(22) xor crc_i(5) xor crc_i(3) xor crc_data_in(19) xor crc_i(19) xor crc_i(2) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(14) xor crc_data_in(18) xor crc_i(18) xor crc_i(14) xor crc_data_in(7) xor crc_data_in(10) xor crc_data_in(25) xor crc_i(1) xor crc_i(25) xor crc_i(10) xor crc_data_in(13) xor crc_data_in(31) xor crc_i(7) xor crc_i(31) xor crc_i(13);
crc_c(14) <= crc_data_in(2) xor crc_data_in(3) xor crc_data_in(4) xor crc_data_in(6) xor crc_data_in(7) xor crc_data_in(17) xor crc_i(7) xor crc_i(17) xor crc_data_in(23) xor crc_i(23) xor crc_i(6) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_i(3) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(15) xor crc_data_in(19) xor crc_i(19) xor crc_i(15) xor crc_data_in(8) xor crc_data_in(11) xor crc_data_in(26) xor crc_i(2) xor crc_i(26) xor crc_i(11) xor crc_data_in(14) xor crc_i(8) xor crc_i(14);
crc_c(15) <= crc_data_in(3) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(7) xor crc_data_in(8) xor crc_data_in(18) xor crc_i(8) xor crc_i(18) xor crc_data_in(24) xor crc_i(24) xor crc_i(7) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_i(4) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(16) xor crc_data_in(20) xor crc_i(20) xor crc_i(16) xor crc_data_in(9) xor crc_data_in(12) xor crc_data_in(27) xor crc_i(3) xor crc_i(27) xor crc_i(12) xor crc_data_in(15) xor crc_i(9) xor crc_i(15);
crc_c(16) <= crc_data_in(0) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(8) xor crc_data_in(19) xor crc_i(19) xor crc_i(8) xor crc_data_in(22) xor crc_i(22) xor crc_i(5) xor crc_data_in(17) xor crc_data_in(21) xor crc_i(21) xor crc_i(17) xor crc_data_in(13) xor crc_i(4) xor crc_i(13) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(26) xor crc_i(26) xor crc_data_in(12) xor crc_data_in(30) xor crc_i(30) xor crc_i(12);
crc_c(17) <= crc_data_in(1) xor crc_data_in(5) xor crc_data_in(6) xor crc_data_in(9) xor crc_data_in(20) xor crc_i(20) xor crc_i(9) xor crc_data_in(23) xor crc_i(23) xor crc_i(6) xor crc_data_in(18) xor crc_data_in(22) xor crc_i(22) xor crc_i(18) xor crc_data_in(14) xor crc_i(5) xor crc_i(14) xor crc_data_in(25) xor crc_i(1) xor crc_i(25) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(13) xor crc_data_in(31) xor crc_i(31) xor crc_i(13);
crc_c(18) <= crc_data_in(2) xor crc_data_in(6) xor crc_data_in(7) xor crc_data_in(10) xor crc_data_in(21) xor crc_i(21) xor crc_i(10) xor crc_data_in(24) xor crc_i(24) xor crc_i(7) xor crc_data_in(19) xor crc_data_in(23) xor crc_i(23) xor crc_i(19) xor crc_data_in(15) xor crc_i(6) xor crc_i(15) xor crc_data_in(26) xor crc_i(2) xor crc_i(26) xor crc_data_in(31) xor crc_i(31) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(14) xor crc_i(14);
crc_c(19) <= crc_data_in(3) xor crc_data_in(7) xor crc_data_in(8) xor crc_data_in(11) xor crc_data_in(22) xor crc_i(22) xor crc_i(11) xor crc_data_in(25) xor crc_i(25) xor crc_i(8) xor crc_data_in(20) xor crc_data_in(24) xor crc_i(24) xor crc_i(20) xor crc_data_in(16) xor crc_i(7) xor crc_i(16) xor crc_data_in(27) xor crc_i(3) xor crc_i(27) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(15) xor crc_i(15);
crc_c(20) <= crc_data_in(4) xor crc_data_in(8) xor crc_data_in(9) xor crc_data_in(12) xor crc_data_in(23) xor crc_i(23) xor crc_i(12) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(21) xor crc_data_in(25) xor crc_i(25) xor crc_i(21) xor crc_data_in(17) xor crc_i(8) xor crc_i(17) xor crc_data_in(28) xor crc_i(4) xor crc_i(28) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(16) xor crc_i(16);
crc_c(21) <= crc_data_in(5) xor crc_data_in(9) xor crc_data_in(10) xor crc_data_in(13) xor crc_data_in(24) xor crc_i(24) xor crc_i(13) xor crc_data_in(27) xor crc_i(27) xor crc_i(10) xor crc_data_in(22) xor crc_data_in(26) xor crc_i(26) xor crc_i(22) xor crc_data_in(18) xor crc_i(9) xor crc_i(18) xor crc_data_in(29) xor crc_i(5) xor crc_i(29) xor crc_data_in(31) xor crc_i(31) xor crc_data_in(17) xor crc_i(17);
crc_c(22) <= crc_data_in(0) xor crc_data_in(11) xor crc_data_in(14) xor crc_i(14) xor crc_i(11) xor crc_data_in(23) xor crc_data_in(27) xor crc_i(27) xor crc_i(23) xor crc_data_in(19) xor crc_i(19) xor crc_data_in(18) xor crc_i(18) xor crc_data_in(9) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(12) xor crc_data_in(16) xor crc_i(16) xor crc_data_in(31) xor crc_i(31) xor crc_i(12);
crc_c(23) <= crc_data_in(0) xor crc_data_in(1) xor crc_data_in(15) xor crc_i(15) xor crc_data_in(20) xor crc_i(20) xor crc_data_in(19) xor crc_i(19) xor crc_i(1) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(13) xor crc_data_in(17) xor crc_i(17) xor crc_i(13) xor crc_data_in(6) xor crc_data_in(9) xor crc_i(0) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(26) xor crc_i(26) xor crc_i(9) xor crc_data_in(16) xor crc_i(6) xor crc_i(16) xor crc_data_in(31) xor crc_i(31);
crc_c(24) <= crc_data_in(1) xor crc_data_in(2) xor crc_data_in(16) xor crc_i(16) xor crc_data_in(21) xor crc_i(21) xor crc_data_in(20) xor crc_i(20) xor crc_i(2) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(14) xor crc_data_in(18) xor crc_i(18) xor crc_i(14) xor crc_data_in(7) xor crc_data_in(10) xor crc_i(1) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(27) xor crc_i(27) xor crc_i(10) xor crc_data_in(17) xor crc_i(7) xor crc_i(17);
crc_c(25) <= crc_data_in(2) xor crc_data_in(3) xor crc_data_in(17) xor crc_i(17) xor crc_data_in(22) xor crc_i(22) xor crc_data_in(21) xor crc_i(21) xor crc_i(3) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(15) xor crc_data_in(19) xor crc_i(19) xor crc_i(15) xor crc_data_in(8) xor crc_data_in(11) xor crc_i(2) xor crc_data_in(31) xor crc_i(31) xor crc_data_in(28) xor crc_i(28) xor crc_i(11) xor crc_data_in(18) xor crc_i(8) xor crc_i(18);
crc_c(26) <= crc_data_in(0) xor crc_data_in(3) xor crc_data_in(4) xor crc_data_in(18) xor crc_i(18) xor crc_data_in(23) xor crc_i(23) xor crc_data_in(22) xor crc_i(22) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_i(3) xor crc_data_in(19) xor crc_i(19) xor crc_data_in(6) xor crc_data_in(10) xor crc_data_in(24) xor crc_i(0) xor crc_i(24) xor crc_data_in(28) xor crc_i(28) xor crc_i(10) xor crc_data_in(26) xor crc_i(26) xor crc_data_in(25) xor crc_i(25) xor crc_i(6) xor crc_data_in(31) xor crc_i(31);
crc_c(27) <= crc_data_in(1) xor crc_data_in(4) xor crc_data_in(5) xor crc_data_in(19) xor crc_i(19) xor crc_data_in(24) xor crc_i(24) xor crc_data_in(23) xor crc_i(23) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_i(4) xor crc_data_in(20) xor crc_i(20) xor crc_data_in(7) xor crc_data_in(11) xor crc_data_in(25) xor crc_i(1) xor crc_i(25) xor crc_data_in(29) xor crc_i(29) xor crc_i(11) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(26) xor crc_i(26) xor crc_i(7);
crc_c(28) <= crc_data_in(2) xor crc_data_in(5) xor crc_data_in(6) xor crc_data_in(20) xor crc_i(20) xor crc_data_in(25) xor crc_i(25) xor crc_data_in(24) xor crc_i(24) xor crc_i(6) xor crc_data_in(22) xor crc_i(22) xor crc_i(5) xor crc_data_in(21) xor crc_i(21) xor crc_data_in(8) xor crc_data_in(12) xor crc_data_in(26) xor crc_i(2) xor crc_i(26) xor crc_data_in(30) xor crc_i(30) xor crc_i(12) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(27) xor crc_i(27) xor crc_i(8);
crc_c(29) <= crc_data_in(3) xor crc_data_in(6) xor crc_data_in(7) xor crc_data_in(21) xor crc_i(21) xor crc_data_in(26) xor crc_i(26) xor crc_data_in(25) xor crc_i(25) xor crc_i(7) xor crc_data_in(23) xor crc_i(23) xor crc_i(6) xor crc_data_in(22) xor crc_i(22) xor crc_data_in(9) xor crc_data_in(13) xor crc_data_in(27) xor crc_i(3) xor crc_i(27) xor crc_data_in(31) xor crc_i(31) xor crc_i(13) xor crc_data_in(29) xor crc_i(29) xor crc_data_in(28) xor crc_i(28) xor crc_i(9);
crc_c(30) <= crc_data_in(4) xor crc_data_in(7) xor crc_data_in(8) xor crc_data_in(22) xor crc_i(22) xor crc_data_in(27) xor crc_i(27) xor crc_data_in(26) xor crc_i(26) xor crc_i(8) xor crc_data_in(24) xor crc_i(24) xor crc_i(7) xor crc_data_in(23) xor crc_i(23) xor crc_data_in(10) xor crc_data_in(14) xor crc_data_in(28) xor crc_i(4) xor crc_i(28) xor crc_i(14) xor crc_data_in(30) xor crc_i(30) xor crc_data_in(29) xor crc_i(29) xor crc_i(10);
crc_c(31) <= crc_data_in(5) xor crc_data_in(8) xor crc_data_in(9) xor crc_data_in(23) xor crc_i(23) xor crc_data_in(28) xor crc_i(28) xor crc_data_in(27) xor crc_i(27) xor crc_i(9) xor crc_data_in(25) xor crc_i(25) xor crc_i(8) xor crc_data_in(24) xor crc_i(24) xor crc_data_in(11) xor crc_data_in(15) xor crc_data_in(29) xor crc_i(5) xor crc_i(29) xor crc_i(15) xor crc_data_in(31) xor crc_i(31) xor crc_data_in(30) xor crc_i(30) xor crc_i(11);

crc_gen_process : process(clk, rst_n)
begin
 if(rst_n = '0') then
    crc_r <= crc_const;				-- reset the valid calculated crc to be the seed
 elsif(rising_edge(clk)) then
    if(crc_data_valid = '1') then
         crc_r <= crc_c;			-- if the input data are valid, save the calculated crc
    end if;
 end if;
end process crc_gen_process;

crc_out <= crc_r;					-- assign the output to be the valid calculated crc

end behave;